module PresentpLayer(
	input wire [63:0] inData,
	output wire [63:0] outData
);

assign outData[0] = inData[0];
assign outData[16] = inData[1];
assign outData[32] = inData[2];
assign outData[48] = inData[3];
assign outData[1] = inData[4];
assign outData[17] = inData[5];
assign outData[33] = inData[6];
assign outData[49] = inData[7];
assign outData[2] = inData[8];
assign outData[18] = inData[9];
assign outData[34] = inData[10];
assign outData[50] = inData[11];
assign outData[3] = inData[12];
assign outData[19] = inData[13];
assign outData[35] = inData[14];
assign outData[51] = inData[15];
assign outData[4] = inData[16];
assign outData[20] = inData[17];
assign outData[36] = inData[18];
assign outData[52] = inData[19];
assign outData[5] = inData[20];
assign outData[21] = inData[21];
assign outData[37] = inData[22];
assign outData[53] = inData[23];
assign outData[6] = inData[24];
assign outData[22] = inData[25];
assign outData[38] = inData[26];
assign outData[54] = inData[27];
assign outData[7] = inData[28];
assign outData[23] = inData[29];
assign outData[39] = inData[30];
assign outData[55] = inData[31];
assign outData[8] = inData[32];
assign outData[24] = inData[33];
assign outData[40] = inData[34];
assign outData[56] = inData[35];
assign outData[9] = inData[36];
assign outData[25] = inData[37];
assign outData[41] = inData[38];
assign outData[57] = inData[39];
assign outData[10] = inData[40];
assign outData[26] = inData[41];
assign outData[42] = inData[42];
assign outData[58] = inData[43];
assign outData[11] = inData[44];
assign outData[27] = inData[45];
assign outData[43] = inData[46];
assign outData[59] = inData[47];
assign outData[12] = inData[48];
assign outData[28] = inData[49];
assign outData[44] = inData[50];
assign outData[60] = inData[51];
assign outData[13] = inData[52];
assign outData[29] = inData[53];
assign outData[45] = inData[54];
assign outData[61] = inData[55];
assign outData[14] = inData[56];
assign outData[30] = inData[57];
assign outData[46] = inData[58];
assign outData[62] = inData[59];
assign outData[15] = inData[60];
assign outData[31] = inData[61];
assign outData[47] = inData[62];
assign outData[63] = inData[63];
endmodule 